//What happens when an enum variable is assigned with the last valid value and the next method is used to do the next assignment?

answer : when the value is already a last valid  but u call next then it show the (x) unknown
