//Why can’t we use a foreach loop for popping all the elements in a queue?  

For each is read only modify panna kudathu 

Pop panna queue size change aagum, so for each confuse agum and it  lead to an error 

Instead we can use the while loop
